class derived_test0 extends abstract_test;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction


  `uvm_component_utils(derived_test0)

endclass
