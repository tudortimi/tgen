module top;

  import tests::*;

  initial
    uvm_pkg::run_test();

endmodule
