package tests;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "sequence0.svh"
  `include "sequence1.svh"

  `include "test0.svh"
  `include "test1.svh"

  `include "abstract_test.svh"
  `include "derived_test0.svh"
  `include "derived_test1.svh"

endpackage
